module ALU(
    input [7:0]A,
    input [7:0]B,
    input [2:0]op,
    output reg [7:0]S //??always???reg???
);
    always@(*)//?????????????
    begin
      case(op)
        3'b000:S = A + B; //?op?000???
        3'b001:S = A - B; //?op?001???
        default:S = 8'bx; //?op????????
      endcase
    end  
endmodule
