library verilog;
use verilog.vl_types.all;
entity test_FSM_counter is
end test_FSM_counter;
