library verilog;
use verilog.vl_types.all;
entity RYG_FSM_test is
end RYG_FSM_test;
