library verilog;
use verilog.vl_types.all;
entity CounterWithController_test is
end CounterWithController_test;
