library verilog;
use verilog.vl_types.all;
entity test_pipeline_ALU is
end test_pipeline_ALU;
