module test_clock;
  reg clk, reset;
  clock clock1(
    .clk(clk),
    .reset(reset)
  );

always #5 clk = ~clk;//?5????clk???

initial
  begin
    clk = 0;reset = 1;//?????
    #10 reset = 0;//10?????????
    #25000 $stop;//25000???????
  end
endmodule
