library verilog;
use verilog.vl_types.all;
entity test_clock is
end test_clock;
