library verilog;
use verilog.vl_types.all;
entity test_BCD_counter is
end test_BCD_counter;
